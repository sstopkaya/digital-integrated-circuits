* SPICE3 file created from AOI22.ext - technology: scmos

M1000 Vdd A a_n27_n9# Vdd pmos w=6u l=2u
+  ad=48p pd=28u as=120p ps=76u
M1001 a_n27_n9# B Vdd Vdd pmos w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y C a_n27_n9# Vdd pmos w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1003 a_n27_n9# D Y Vdd pmos w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_n19_n33# A GND Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=60p ps=44u
M1005 Y B a_n19_n33# Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1006 a_1_n33# C Y Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1007 GND D a_1_n33# Gnd nmos w=5u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Y gnd! 7.4fF
C1 Vdd gnd! 10.7fF
C2 a_n27_n9# gnd! 11.8fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    B     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin2    C     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin3    D     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
