magic
tech scmos
timestamp 1605730781
<< polysilicon >>
rect -15 10 -13 12
rect -7 10 -5 12
rect 1 10 3 12
rect -15 -18 -13 7
rect -7 -11 -5 7
rect 1 -4 3 7
rect -15 -25 -13 -22
rect -7 -25 -5 -15
rect 1 -25 3 -8
rect -15 -30 -13 -28
rect -7 -30 -5 -28
rect 1 -30 3 -28
<< ndiffusion >>
rect -16 -28 -15 -25
rect -13 -28 -7 -25
rect -5 -28 1 -25
rect 3 -28 6 -25
<< pdiffusion >>
rect -16 7 -15 10
rect -13 7 -12 10
rect -8 7 -7 10
rect -5 7 -4 10
rect 0 7 1 10
rect 3 7 6 10
<< metal1 >>
rect -20 14 -8 18
rect -4 14 12 18
rect -20 10 -16 14
rect -4 10 0 14
rect -12 3 -8 6
rect 6 3 10 6
rect -12 -1 10 3
rect -20 -8 -1 -4
rect 6 -11 10 -1
rect -20 -15 -9 -11
rect 6 -15 12 -11
rect -20 -22 -17 -18
rect 6 -24 10 -15
rect -20 -32 -16 -29
rect -20 -36 -8 -32
rect -4 -36 10 -32
<< ntransistor >>
rect -15 -28 -13 -25
rect -7 -28 -5 -25
rect 1 -28 3 -25
<< ptransistor >>
rect -15 7 -13 10
rect -7 7 -5 10
rect 1 7 3 10
<< polycontact >>
rect -1 -8 3 -4
rect -9 -15 -5 -11
rect -17 -22 -13 -18
<< ndcontact >>
rect -20 -29 -16 -25
rect 6 -28 10 -24
<< pdcontact >>
rect -20 6 -16 10
rect -12 6 -8 10
rect -4 6 0 10
rect 6 6 10 10
<< psubstratepcontact >>
rect -8 -36 -4 -32
<< nsubstratencontact >>
rect -8 14 -4 18
<< labels >>
rlabel metal1 11 16 11 18 6 Vdd
rlabel metal1 -19 -7 -19 -5 3 A
rlabel metal1 -19 -14 -19 -12 3 B
rlabel metal1 -19 -21 -19 -19 3 C
rlabel metal1 11 -14 11 -12 7 Y
rlabel metal1 7 -36 7 -34 8 GND
<< end >>
