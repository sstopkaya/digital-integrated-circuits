* SPICE3 file created from NAND3.ext - technology: scmos

M1000 Y C Vdd Vdd pmos w=3u l=2u
+  ad=47p pd=42u as=41p ps=38u
M1001 Vdd B Y Vdd pmos w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A Vdd Vdd pmos w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_n13_n28# C GND Gnd nmos w=3u l=2u
+  ad=18p pd=18u as=19p ps=18u
M1004 a_n5_n28# B a_n13_n28# Gnd nmos w=3u l=2u
+  ad=18p pd=18u as=0p ps=0u
M1005 Y A a_n5_n28# Gnd nmos w=3u l=2u
+  ad=25p pd=22u as=0p ps=0u
C0 Y gnd! 9.7fF
C1 Vdd gnd! 6.8fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    B     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin2    C     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
