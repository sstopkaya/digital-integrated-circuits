magic
tech scmos
timestamp 1605714479
<< polysilicon >>
rect 0 20 2 23
rect 0 12 2 16
rect -4 10 2 12
rect 0 6 2 10
rect 0 0 2 2
<< ndiffusion >>
rect -1 2 0 6
rect 2 2 3 6
<< pdiffusion >>
rect -1 16 0 20
rect 2 16 3 20
<< metal1 >>
rect -11 24 -9 28
rect -5 20 -1 28
rect 3 24 7 28
rect 11 24 14 28
rect 3 13 7 16
rect -10 9 -8 13
rect 3 9 11 13
rect 3 6 7 9
rect -5 -6 -1 2
rect 3 -6 7 -2
rect 11 -6 14 -2
<< ntransistor >>
rect 0 2 2 6
<< ptransistor >>
rect 0 16 2 20
<< polycontact >>
rect -8 9 -4 13
<< ndcontact >>
rect -5 2 -1 6
rect 3 2 7 6
<< pdcontact >>
rect -5 16 -1 20
rect 3 16 7 20
<< psubstratepcontact >>
rect -9 -6 -5 -2
rect -1 -6 3 -2
rect 7 -6 11 -2
<< nsubstratencontact >>
rect -9 24 -5 28
rect -1 24 3 28
rect 7 24 11 28
<< labels >>
rlabel metal1 11 11 11 13 7 Y
rlabel metal1 14 -6 14 -4 8 GND
rlabel metal1 14 26 14 28 6 Vdd
rlabel metal1 -10 11 -10 13 3 A
<< end >>
