* SPICE3 file created from MUX2x1.ext - technology: scmos

M1000 Vdd D0 a_n27_n9# Vdd pmos w=6u l=2u
+  ad=48p pd=28u as=120p ps=76u
M1001 a_n27_n9# Sn Vdd Vdd pmos w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y S a_n27_n9# Vdd pmos w=6u l=2u
+  ad=48p pd=28u as=0p ps=0u
M1003 a_n27_n9# D1 Y Vdd pmos w=6u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_n19_n33# D0 GND Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=60p ps=44u
M1005 Y Sn a_n19_n33# Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1006 a_1_n33# S Y Gnd nmos w=5u l=2u
+  ad=40p pd=26u as=0p ps=0u
M1007 GND D1 a_1_n33# Gnd nmos w=5u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Y gnd! 7.2fF
C1 a_n27_n9# gnd! 11.5fF
C2 S gnd! 6.4fF
C3 Sn gnd! 6.4fF
C4 Vdd gnd! 8.5fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     D0     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    Sn     GND    PWL(   0   2.5    4N  2.5    4.1N 0   8N  0  8.1N  2.5  ) 
Vin2    S      GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin3    D1     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
