magic
tech scmos
timestamp 1605752816
<< polysilicon >>
rect -28 1 -26 4
rect -20 1 -18 4
rect -8 1 -6 4
rect 0 1 2 4
rect -28 -25 -26 -6
rect -20 -25 -18 -6
rect -8 -25 -6 -6
rect 0 -25 2 -6
rect -28 -31 -26 -29
rect -20 -31 -18 -29
rect -8 -31 -6 -29
rect 0 -31 2 -29
<< ndiffusion >>
rect -29 -29 -28 -25
rect -26 -29 -25 -25
rect -21 -29 -20 -25
rect -18 -29 -15 -25
rect -11 -29 -8 -25
rect -6 -29 -5 -25
rect -1 -29 0 -25
rect 2 -29 3 -25
<< pdiffusion >>
rect -29 -6 -28 1
rect -26 -6 -20 1
rect -18 -6 -15 1
rect -11 -6 -8 1
rect -6 -6 0 1
rect 2 -6 3 1
<< metal1 >>
rect -33 7 -25 11
rect -21 7 -15 11
rect -11 7 -4 11
rect 0 7 7 11
rect -33 6 7 7
rect -33 1 -29 6
rect 3 1 7 6
rect -15 -11 -11 -6
rect -15 -15 9 -11
rect -33 -22 -11 -18
rect -33 -25 -29 -22
rect -15 -25 -11 -22
rect -25 -40 -21 -29
rect -5 -25 -1 -15
rect -15 -33 -11 -29
rect 3 -33 7 -29
rect -15 -37 7 -33
rect -33 -41 9 -40
rect -33 -45 -25 -41
rect -21 -45 -14 -41
rect -10 -45 -3 -41
rect 1 -45 9 -41
<< ntransistor >>
rect -28 -29 -26 -25
rect -20 -29 -18 -25
rect -8 -29 -6 -25
rect 0 -29 2 -25
<< ptransistor >>
rect -28 -6 -26 1
rect -20 -6 -18 1
rect -8 -6 -6 1
rect 0 -6 2 1
<< ndcontact >>
rect -33 -29 -29 -25
rect -25 -29 -21 -25
rect -15 -29 -11 -25
rect -5 -29 -1 -25
rect 3 -29 7 -25
<< pdcontact >>
rect -33 -6 -29 1
rect -15 -6 -11 1
rect 3 -6 7 1
<< psubstratepcontact >>
rect -25 -45 -21 -41
rect -14 -45 -10 -41
rect -3 -45 1 -41
<< nsubstratencontact >>
rect -25 7 -21 11
rect -15 7 -11 11
rect -4 7 0 11
<< labels >>
rlabel polysilicon -20 4 -18 4 1 B
rlabel polysilicon -28 4 -26 4 1 A
rlabel metal1 5 -43 5 -41 1 GND
rlabel polysilicon -8 4 -6 4 1 C
rlabel polysilicon 0 4 2 4 1 D
rlabel metal1 4 10 5 10 6 Vdd
rlabel metal1 6 -14 6 -12 7 Y
<< end >>
