* SPICE3 file created from NOR2.ext - technology: scmos

M1000 a_n22_0# B Vdd Vdd pmos w=3u l=2u
+  ad=24p pd=22u as=19p ps=18u
M1001 Y A a_n22_0# Vdd pmos w=3u l=2u
+  ad=22p pd=20u as=0p ps=0u
M1002 Y B GND Gnd nmos w=3u l=2u
+  ad=28p pd=24u as=38p ps=36u
M1003 GND A Y Gnd nmos w=3u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Y gnd! 5.3fF
C1 Vdd gnd! 3.6fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    B     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
