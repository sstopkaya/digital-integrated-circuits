magic
tech scmos
timestamp 1605749306
<< polysilicon >>
rect -21 -3 -19 -1
rect -11 -3 -9 -1
rect -1 -3 1 -1
rect 9 -3 11 -1
rect -21 -28 -19 -9
rect -11 -28 -9 -9
rect -1 -28 1 -9
rect 9 -28 11 -9
rect -21 -35 -19 -33
rect -11 -35 -9 -33
rect -1 -35 1 -33
rect 9 -35 11 -33
<< ndiffusion >>
rect -23 -33 -21 -28
rect -19 -33 -11 -28
rect -9 -33 -7 -28
rect -3 -33 -1 -28
rect 1 -33 9 -28
rect 11 -33 13 -28
<< pdiffusion >>
rect -23 -9 -21 -3
rect -19 -9 -17 -3
rect -13 -9 -11 -3
rect -9 -9 -7 -3
rect -3 -9 -1 -3
rect 1 -9 3 -3
rect 7 -9 9 -3
rect 11 -9 13 -3
<< metal1 >>
rect -27 8 19 12
rect -17 -3 -13 8
rect -7 1 17 5
rect -7 -3 -3 1
rect 13 -3 17 1
rect -27 -13 -23 -9
rect -7 -13 -3 -9
rect -27 -17 -3 -13
rect 3 -20 7 -9
rect -7 -24 19 -20
rect -7 -28 -3 -24
rect -27 -37 -23 -33
rect 13 -37 17 -33
rect -27 -41 19 -37
<< ntransistor >>
rect -21 -33 -19 -28
rect -11 -33 -9 -28
rect -1 -33 1 -28
rect 9 -33 11 -28
<< ptransistor >>
rect -21 -9 -19 -3
rect -11 -9 -9 -3
rect -1 -9 1 -3
rect 9 -9 11 -3
<< ndcontact >>
rect -27 -33 -23 -28
rect -7 -33 -3 -28
rect 13 -33 17 -28
<< pdcontact >>
rect -27 -9 -23 -3
rect -17 -9 -13 -3
rect -7 -9 -3 -3
rect 3 -9 7 -3
rect 13 -9 17 -3
<< labels >>
rlabel metal1 17 -23 17 -21 7 Y
rlabel metal1 17 -40 17 -38 8 GND
rlabel metal1 16 10 16 12 6 Vdd
rlabel polysilicon -21 -1 -19 -1 1 A
rlabel polysilicon -11 -1 -9 -1 1 B
rlabel polysilicon -1 -1 1 -1 1 C
rlabel polysilicon 9 -1 11 -1 1 D
<< end >>
