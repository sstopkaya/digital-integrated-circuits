magic
tech scmos
timestamp 1605744964
<< polysilicon >>
rect -28 1 -26 4
rect -20 1 -18 4
rect -7 1 -5 4
rect 1 1 3 4
rect -28 -25 -26 -6
rect -20 -25 -18 -6
rect -7 -25 -5 -6
rect 1 -25 3 -6
rect -28 -31 -26 -29
rect -20 -31 -18 -29
rect -7 -31 -5 -29
rect 1 -31 3 -29
<< ndiffusion >>
rect -29 -29 -28 -25
rect -26 -29 -25 -25
rect -21 -29 -20 -25
rect -18 -29 -15 -25
rect -11 -29 -7 -25
rect -5 -29 -4 -25
rect 0 -29 1 -25
rect 3 -29 4 -25
<< pdiffusion >>
rect -29 -6 -28 1
rect -26 -6 -20 1
rect -18 -6 -15 1
rect -11 -6 -7 1
rect -5 -6 1 1
rect 3 -6 4 1
<< metal1 >>
rect -31 7 -25 11
rect -21 7 -15 11
rect -11 7 -4 11
rect 0 7 5 11
rect -31 6 5 7
rect -15 1 -11 6
rect -33 -10 -29 -6
rect 4 -10 8 -6
rect -33 -14 10 -10
rect -25 -25 -21 -14
rect -15 -22 8 -18
rect -15 -25 -11 -22
rect 4 -25 8 -22
rect -33 -33 -29 -29
rect -15 -33 -11 -29
rect -33 -37 -11 -33
rect -4 -40 0 -29
rect -33 -41 8 -40
rect -33 -45 -26 -41
rect -22 -45 -15 -41
rect -11 -45 -4 -41
rect 0 -45 8 -41
<< ntransistor >>
rect -28 -29 -26 -25
rect -20 -29 -18 -25
rect -7 -29 -5 -25
rect 1 -29 3 -25
<< ptransistor >>
rect -28 -6 -26 1
rect -20 -6 -18 1
rect -7 -6 -5 1
rect 1 -6 3 1
<< ndcontact >>
rect -33 -29 -29 -25
rect -25 -29 -21 -25
rect -15 -29 -11 -25
rect -4 -29 0 -25
rect 4 -29 8 -25
<< pdcontact >>
rect -33 -6 -29 1
rect -15 -6 -11 1
rect 4 -6 8 1
<< psubstratepcontact >>
rect -26 -45 -22 -41
rect -15 -45 -11 -41
rect -4 -45 0 -41
<< nsubstratencontact >>
rect -25 7 -21 11
rect -15 7 -11 11
rect -4 7 0 11
<< labels >>
rlabel polysilicon -20 4 -18 4 1 B
rlabel polysilicon -7 4 -5 4 1 A
rlabel polysilicon 1 4 3 4 1 Bn
rlabel metal1 8 -13 8 -11 7 Y
rlabel polysilicon -28 4 -26 4 1 An
rlabel metal1 4 -43 4 -41 1 GND
rlabel metal1 2 10 3 10 5 Vdd
<< end >>
