* SPICE3 file created from INV.ext - technology: scmos

M1000 Y A Vdd Vdd pmos w=4u l=2u
+  ad=20p pd=18u as=20p ps=18u
M1001 Y A GND Gnd nmos w=4u l=2u
+  ad=20p pd=18u as=20p ps=18u
C0 Y gnd! 2.6fF
C1 Vdd gnd! 3.2fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    4N  2.5    4.1N 0   8N  0  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END

