* SPICE3 file created from XNOR2.ext - technology: scmos

M1000 a_n26_n6# A Y Vdd pmos w=7u l=2u
+  ad=42p pd=26u as=70p ps=48u
M1001 Vdd B a_n26_n6# Vdd pmos w=7u l=2u
+  ad=77p pd=36u as=0p ps=0u
M1002 a_n5_n6# An Vdd Vdd pmos w=7u l=2u
+  ad=42p pd=26u as=0p ps=0u
M1003 Y Bn a_n5_n6# Vdd pmos w=7u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A a_n33_n29# Gnd nmos w=4u l=2u
+  ad=24p pd=20u as=84p ps=66u
M1005 a_n33_n29# B Y Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1006 GND An a_n33_n29# Gnd nmos w=4u l=2u
+  ad=24p pd=20u as=0p ps=0u
M1007 a_n33_n29# Bn GND Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 a_n33_n29# gnd! 10.8fF
C1 Y gnd! 11.1fF
C2 Vdd gnd! 7.1fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A      GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    B      GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin2    An     GND    PWL(   0   2.5    4N  2.5    4.1N 0   8N  0  8.1N  2.5  ) 
Vin3    Bn     GND    PWL(   0   2.5    4N  2.5    4.1N 0   8N  0  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
