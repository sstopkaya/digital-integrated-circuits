* SPICE3 file created from NOR3.ext - technology: scmos

M1000 a_n7_1# C Vdd Vdd pmos w=6u l=2u
+  ad=12p pd=16u as=30p ps=22u
M1001 a_n3_1# B a_n7_1# Vdd pmos w=6u l=2u
+  ad=12p pd=16u as=0p ps=0u
M1002 Y A a_n3_1# Vdd pmos w=6u l=2u
+  ad=30p pd=22u as=0p ps=0u
M1003 Y C GND Gnd nmos w=4u l=2u
+  ad=44p pd=38u as=44p ps=38u
M1004 GND B Y Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A GND Gnd nmos w=4u l=2u
+  ad=0p pd=0u as=0p ps=0u
C0 Y gnd! 11.4fF
C1 Vdd gnd! 7.0fF

VCC    VDD     GND     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3    T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --    --  --  ---- -- 
Vin     A     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin1    B     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 
Vin2    C     GND    PWL(   0   2.5    4N  2.5    4.1N 2.5   8N  2.5  8.1N  2.5  ) 


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1


* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
